LIBRARY ieee;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_1164.ALL;

ENTITY ordBits IS
	PORT(ordIn: IN unsigned (4 DOWNTO 0);
		  ordOut: OUT unsigned(15 DOWNTO 0));
END ENTITY;


ARCHITECTURE ordBits OF ordBits IS

BEGIN
	ordOut <= "0000000000000000" WHEN ordIn = "00000" ELSE
				 "1000000000000000" WHEN ordIn = "00001" ELSE
				 "1100000000000000" WHEN ordIn = "00010" ELSE
				 "1110000000000000" WHEN ordIn = "00011" ELSE
				 "1111000000000000" WHEN ordIn = "00100" ELSE
				 "1111100000000000" WHEN ordIn = "00101" ELSE
				 "1111110000000000" WHEN ordIn = "00110" ELSE
				 "1111111000000000" WHEN ordIn = "00111" ELSE
				 "1111111100000000" WHEN ordIn = "01000" ELSE
				 "1111111110000000" WHEN ordIn = "01001" ELSE
				 "1111111111000000" WHEN ordIn = "01010" ELSE
				 "1111111111100000" WHEN ordIn = "01011" ELSE
				 "1111111111110000" WHEN ordIn = "01100" ELSE
				 "1111111111111000" WHEN ordIn = "01101" ELSE
				 "1111111111111100" WHEN ordIn = "01110" ELSE
				 "1111111111111110" WHEN ordIn = "01111" ELSE
				 "1111111111111111" WHEN ordIn = "10000" ELSE
				 "XXXXXXXXXXXXXXXX";
END ARCHITECTURE;