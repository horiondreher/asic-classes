LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY Dec_To_Frac IS
	PORT(	DecIn: IN unsigned(3 DOWNTO 0);
			DecOut: OUT unsigned(51 DOWNTO 0));
END ENTITY;

ARCHITECTURE Dec_To_Frac OF Dec_To_Frac IS

TYPE mem IS ARRAY(0 TO 9) OF unsigned(51 DOWNTO 0);
SIGNAL aux: mem := (	"0000000000000000000000000000000000000000000000000000",
							"0001100110011001100110011001100110011001100110011001",
							"0011001100110011001100110011001100110011001100110011",
							"0100110011001100110011001100110011001100110011001100",
							"0110011001100110011001100110011001100110011001100110",
							"1000000000000000000000000000000000000000000000000000",
							"1001100110011001100110011001100110011001100110011001",
							"1011001100110011001100110011001100110011001100110011",
							"1100110011001100110011001100110011001100110011001100",
							"1110011001100110011001100110011001100110011001100110");
SIGNAL address : integer RANGE 0 TO 9 := to_integer(DecIn);					
	
BEGIN

	DecOut <= aux(address);	
	
END ARCHITECTURE;