LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY Cent_To_Frac IS
	PORT(	CentIn: IN unsigned(3 DOWNTO 0);
			CentOut: OUT unsigned(51 DOWNTO 0));
END ENTITY;

ARCHITECTURE Cent_To_Frac OF Cent_To_Frac IS

TYPE mem IS ARRAY(0 TO 9) OF unsigned(51 DOWNTO 0);
SIGNAL aux: mem := (	"0000000000000000000000000000000000000000000000000000",
							"0000001010001111010111000010100011110101110000101000",
							"0000010100011110101110000101000111101011100001010001",
							"0000011110101110000101000111101011100001010001111010",
							"0000101000111101011100001010001111010111000010100011",
							"0000110011001100110011001100110011001100110011001100",
							"0000111101011100001010001111010111000010100011110101",
							"0001000111101011100001010001111010111000010100011110",
							"0001010001111010111000010100011110101110000101000111",
							"0001011100001010001111010111000010100011110101110000");
SIGNAL address : integer RANGE 0 TO 9 := to_integer(CentIn);				
	
BEGIN

	CentOut <= aux(address);	
	
END ARCHITECTURE;