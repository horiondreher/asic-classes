LIBRARY ieee;
USE ieee.numeric_std.ALL;

ENTITY inBlock_4bits IS
	PORT(SW : IN unsigned(15 DOWNTO 0); S : OUT unsigned(3 DOWNTO 0));
END ENTITY;

ARCHITECTURE inBlock_4bits OF inBlock_4bits IS
BEGIN 
	WITH SW SELECT
		S <=  "0000" WHEN "0000000000000001",
				"0001" WHEN "0000000000000010",
				"0010" WHEN "0000000000000100",
				"0011" WHEN "0000000000001000",
				"0100" WHEN "0000000000010000",
				"0101" WHEN "0000000000100000",
				"0110" WHEN "0000000001000000",
				"0111" WHEN "0000000010000000",
				"1000" WHEN "0000000100000000",
				"1001" WHEN "0000001000000000",
				"1010" WHEN "0000010000000000",
				"1011" WHEN "0000100000000000",
				"1100" WHEN "0001000000000000",
				"1101" WHEN "0010000000000000",
				"1110" WHEN "0100000000000000",
				"1111" WHEN "1000000000000000",
				"XXXX" WHEN OTHERS;
END ARCHITECTURE;